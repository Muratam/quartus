library verilog;
use verilog.vl_types.all;
entity x16_vlg_tst is
end x16_vlg_tst;
