library verilog;
use verilog.vl_types.all;
entity x16 is
    port(
        x16_o0          : out    vl_logic;
        x16_i0          : in     vl_logic;
        x16_o1          : out    vl_logic;
        x16_i2          : in     vl_logic;
        x16_o2          : out    vl_logic;
        x16_i1          : in     vl_logic;
        x16_o3          : out    vl_logic;
        x16_i3          : in     vl_logic;
        x16_o4          : out    vl_logic;
        x16_o5          : out    vl_logic;
        x16_o6          : out    vl_logic;
        x16_o7          : out    vl_logic
    );
end x16;
